    /**
    * TOP LEVEL MODULE: make_pixel.v
    *  
    * This module is reponsible for drawing all 
    *   
    *
    *
    */


   module make_pixel(
   
        input X_POS,
        input Y_POS,
        input SQ_SIZE,
   
   );
   /**
    * Draws a square of SQ_SIZE to the screen at X_POS and Y_POS
    *
    */

    


   endmodule
