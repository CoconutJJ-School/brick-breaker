
module make_line();
    

endmodule



